`include "width.h"
module tlb
#(
    parameter TLBNUM = 16
)
(
    input  wire                      clk,
    // search port 0 (for fetch)
    input  wire [              18:0] s0_vppn,
    input  wire                      s0_va_bit12,
    input  wire [               9:0] s0_asid,
    output wire                      s0_found,
    output wire [$clog2(TLBNUM)-1:0] s0_index,
    output wire [              19:0] s0_ppn,
    output wire [               5:0] s0_ps,
    output wire [               1:0] s0_plv,
    output wire [               1:0] s0_mat,
    output wire                      s0_d,
    output wire                      s0_v,

    // search port 1 (for load/store)
    input  wire [              18:0] s1_vppn,
    input  wire                      s1_va_bit12,
    input  wire [               9:0] s1_asid,
    output wire                      s1_found,
    output wire [$clog2(TLBNUM)-1:0] s1_index,
    output wire [              19:0] s1_ppn,
    output wire [               5:0] s1_ps,
    output wire [               1:0] s1_plv,
    output wire [               1:0] s1_mat,
    output wire                      s1_d,
    output wire                      s1_v,

    // invtlb opcode
    input  wire                      invtlb_valid,
    input  wire [               4:0] invtlb_op,

    // write port
    input  wire                      we,       //w(rite) e(nable)
    input  wire [$clog2(TLBNUM)-1:0] w_index,
    input  wire                      w_e,
    input  wire [              18:0] w_vppn,
    input  wire [               5:0] w_ps,
    input  wire [               9:0] w_asid,
    input  wire                      w_g,
    input  wire [              19:0] w_ppn0,
    input  wire [               1:0] w_plv0,
    input  wire [               1:0] w_mat0,
    input  wire                      w_d0,
    input  wire                      w_v0,
    input  wire [              19:0] w_ppn1,
    input  wire [               1:0] w_plv1,
    input  wire [               1:0] w_mat1,
    input  wire                      w_d1,
    input  wire                      w_v1,

    // read port
    input  wire [$clog2(TLBNUM)-1:0] r_index,
    output wire                      r_e,
    output wire [              18:0] r_vppn,
    output wire [               5:0] r_ps,
    output wire [               9:0] r_asid,
    output wire                      r_g,
    output wire [              19:0] r_ppn0,
    output wire [               1:0] r_plv0,
    output wire [               1:0] r_mat0,
    output wire                      r_d0,
    output wire                      r_v0,
    output wire [              19:0] r_ppn1,
    output wire [               1:0] r_plv1,
    output wire [               1:0] r_mat1,
    output wire                      r_d1,
    output wire                      r_v1
);
    reg  [TLBNUM-1:0] tlb_e;
    reg  [TLBNUM-1:0] tlb_ps4MB; //pagesize1:4MB,0:4KB
    reg  [      18:0] tlb_vppn   [TLBNUM-1:0];
    reg  [       9:0] tlb_asid   [TLBNUM-1:0];
    reg               tlb_g      [TLBNUM-1:0];
    reg  [      19:0] tlb_ppn0   [TLBNUM-1:0];
    reg  [       1:0] tlb_plv0   [TLBNUM-1:0];
    reg  [       1:0] tlb_mat0   [TLBNUM-1:0];
    reg               tlb_d0     [TLBNUM-1:0];
    reg               tlb_v0     [TLBNUM-1:0];
    reg  [      19:0] tlb_ppn1   [TLBNUM-1:0];
    reg  [       1:0] tlb_plv1   [TLBNUM-1:0];
    reg  [       1:0] tlb_mat1   [TLBNUM-1:0];
    reg               tlb_d1     [TLBNUM-1:0];
    reg               tlb_v1     [TLBNUM-1:0];

    wire [TLBNUM-1:0] match0;
    wire [TLBNUM-1:0] match1;

    wire [TLBNUM-1:0] cond1;
    wire [TLBNUM-1:0] cond2;
    wire [TLBNUM-1:0] cond3;
    wire [TLBNUM-1:0] cond4;

    wire [TLBNUM-1:0] invtlb_mask [31:0];

    genvar i;
    generate
        for (i = 0; i < TLBNUM; i = i + 1) begin
            assign match0[i] = (s0_vppn[18:10] == tlb_vppn[i][18:10])
                                &&(tlb_ps4MB[i] || s0_vppn[9:0] == tlb_vppn[i][9:0])
                                &&((s0_asid == tlb_asid[i]) || tlb_g[i]);
            assign match1[i] = (s1_vppn[18:10] == tlb_vppn[i][18:10])
                                &&(tlb_ps4MB[i] || s1_vppn[9:0] == tlb_vppn[i][9:0])
                                &&((s1_asid == tlb_asid[i]) || tlb_g[i]);
        end    
    endgenerate
    
    generate
        for (i = 0; i < TLBNUM; i = i + 1) begin
            assign cond1[i] = ~tlb_g[i];
            assign cond2[i] = tlb_g[i];
            assign cond3[i] = s1_asid == tlb_asid[i];
            assign cond4[i] = (s1_vppn[18:10] == tlb_vppn[i][18:10]) 
                               && (tlb_ps4MB[i] || s1_vppn[9:0] == tlb_vppn[i][9:0]);
        end
    endgenerate

    assign invtlb_mask[0] = 16'hffff;  
    assign invtlb_mask[1] = 16'hffff;
    assign invtlb_mask[2] = cond2;
    assign invtlb_mask[3] = cond1;
    assign invtlb_mask[4] = cond1 & cond3;
    assign invtlb_mask[5] = cond1 & cond3 & cond4;
    assign invtlb_mask[6] = (cond1 | cond3) & cond4;
    generate
        for (i = 7; i < 32; i = i + 1) begin
            assign invtlb_mask[i] = 16'b0;
        end
    endgenerate


endmodule